`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MrL1Cxn094JIjO1Od2RBtR8jg36cXCYKbrt7DFfFJbN2/N5RBoCdtCQCYIcSp/d
qlTaGHT4srEUdYu3iVhPrrSfKMInILLYRQ+38kBgeBJPp/qR5uNjNV8MOF0LCkJo
lZPqXLvzBi7Y+HpWtSk6AOEBhr9Ss7abOSC2QDiw6xPfvoSN1Ofjbfq7iAVDsNft
7sADiMoQAifXzRbIcBbR9hqXRUoSS7ujJ+qVvf+fuOjB7rOJ3ZqkFrfz+qQ+Ibm4
pNgtRG7oLlTuFRASNcDR9FQLer53oVmcEG9bvb3mSRrnRW2ktGSkkVeiRV6DAn+B
0QKLspv9LL6zhmJSg6L3Obyefdk5zpTr1j+3QGtxTPM7U1efE2gaX4yjTsTmBIcm
cvqgyVZog4OvzZ0OxsQUj36473HDAcM3w9Z2b/8Vvb/UfjdtLK2Ki09fxv1yT7/c
AWZlb+rGmfPa7dgyzQfQLEVzad+Iamb/QnetdIPPS/LitlaMz4atcMCCvdqLkUN9
x2HE8py+qG/xt9rXXXK1a+fDWSDq5ov0MQg8I9IHx0ECeX3pVJFykgeQzttj6ejZ
QifiaRkVg+E7ohVPO9weMUXB8th1GofJkztKMNXgM3WfNerNh6gHSijeZI2m9odN
cKnXGHIOztT1bsXjy9l8Hk0AukeZIZtfbhECQoLmidX1+iPNHK2b5tF2veoaD8Ty
cC/aTYvYlzF0CnXEFUOzlihMVANJsKsE+0KX1WgtxKZV9T3DEylETsoJwOIqvtlr
aZbt0mWMPQwpKm5wk8M5hFQuNO7G8Ix6R6I/D8psGMk/4TgsqOv2GJnA58w2AkIu
JBo52QyZj1hlA+rb472N/e7xaR8qINMNojBFLaaFEC+GQWG3ZUidyhBjmQdf7/4W
1QijVJSJrM75LE2P2zJFjRAa/L1AHIPcTtPjAMHWEH2dB9cp/GeY3/b2qmWHXAvC
RpryJjeO1ZpsDIInOofvx7MiIZCIKyuvTulPP7NjILYGtcs1GGtZPsN2BCF7FxpQ
ys+XVLLg0CN9Us/aJxDat/omkKaI4xSUDiIyjh7/cnOP7UMFgf9Va9CVcNhTeoP0
nfI5rCpfrXR2HiSwbrzGiTpI5ek+76mVjsXdPzHKvixYmDvky99xorCy8NI2sSeo
H3FR2yshhlv0U3oYGTvZA3SWVcBiQQnJViH5nJ040I7/h3w9EEZzQj6ycN9R+IPa
gE+xLUyzsPp/z9ngZxlhg9KR4qPvwHaCTLOYR1cBAZwHX/ORkhIIhN81yJOMVckt
gwOuXwQpwbHzbA/mbzSGrCx7/ihXTDytKGU+qS+XNWtmnejWgZoAh29gtBQ2x7Ez
dwlazuxqH8lvUKEJ3uooqXdb8SQpczFRt81rDr+XpZxRdk1O9nPnuXdPsxi8aLsJ
RQEpfD5iyqlKEg9VwG75lAATv+U21hx2WCHQGNxoESbAIBVSgXWjcNK2htRBpN6G
nV6VCFxtaldgV8L/6LY6fx/dOxA2sDapbYS0GLcjEq5UQySNzwL+Lfcof305TlZB
Ghz/vIM9Tb4GuMT4L8C/j4Y8z62TFj4GlyRnCYhuvqa3bmvM307mlQBN+Nm6Eirq
3whmQlPu//NJtGjsPEvZvEHmsPbuxyHzTVW0Usgd6sck5bORfRqUsCh7W7rKoW6X
/nr9Llrn3lqTVMVsdZjByiG0Si4y8KSUZu6CL8zGeJtGJ/1ScV11wI8gWffUPBQD
r4qwo/NuxNMdg7O+fFaXfBNwldBlRE4Z73w09fW8Wg6ylAp0cD9kD1OxV3RwdcaO
t7GiF08jaQeiqAsE37zIoVBTRypJC0hJzkHapTZnBAMGAHVCVj8EOfZeKRomvnUL
LRd4G3Y0B+/ofs0NLyXwTgcDR0A1uqTuHo1cGrnrpghem1XbVAPbos8sKha3nODd
EFADl9/lyBCeHjU6oNv71MHGTGqB9dcr3n+x8i2dvayw7W56DeE0ZrX04uuBJdsj
KFX3d2G9bx/7R+EoO6v/7hg0N3ccOhXOYpz3VZXFbYVuXGKFoDfYdaDEDMBROfJ1
PmbwNqBbeVgiK7MRY5uxAtXkB+000fOpxZl8E3ITjdTWp5NEnnpLUdktKrRdXXct
MDpfHrHAVxkNnAkL9ITryoYwL9lcpV38PyRmyDNkHT/wGCKLp6YxI74i7A1RokE/
VNXuWB7MtluqTbiMi2I9xnLtP/LA4bScHRR/iIyqFB3Mw85pKU5f8VQNmZzcvC04
mrKWsbYIV1bnK4FEj+fiADp9wbWjfN+eMzNfMv3ApbWmLMCMjUtENNEhKLFqkgUA
4iBNRyidLc5QJlkIOAZ3F4JMKYCrq0+r/Y5C6mN03lg7vNREkk2yGgFpZpOY3RAm
V3R6E3dTJ1HmfAu0CMbaOrSPs4OR0dnKQu14YUSTyMcIXOHdKzZdJqvzoDtEdjrE
mxqSHYlnAS32SNTSkC+V87zdmml4pGSPwcF50Jqn5ouTqNma5EtqXDbXzhTJTeCf
KZpiAslihUX9NFv4balgsDIO/pqw2vx+4lmhZrGshyDCD5HQpEmDKr8Ygwa+05qG
Rt6Hk9rMDf9mw9Rn8l0K3NS12E37p2I3y9eWc6zXdyxsoy7xEzBEUg5ZTMVDAJDe
u1DKp3hx7gyVHSp3uyLyp2vbHHPZdhf08bTrkyENrGMVVXGqeeZU4yE5mM6VY9Ei
KITSO1l5337FX1aX8WjhGKaS6822sDrB6642/DqMD/He/jf7/AgWW7MjINTynDW1
oW89lwjKnK/6mREOQMhelT2V/IYmM9C8AQfW+T5cbnKEvwaaxVdtePkuRKdglXJ8
Vxdvp1924bwG2prGPQmC7gCFvIILSbZgtrT1Ud9DJ9H2O6jIbV8EJUP80jaxuaEE
PXnQcHHc4rsZqXBLXyH/ExsWdkhLIYKMfij+zdlQvzS0/6Fy4SPZKtSEwiyRIIh6
0mweTXHYyBf4LI+pQwNedCa8S0Wtl5J/x3iKrwzdCYXrRmm1M3o6ol1iAWGsMwWK
ka4O292fhhcv5DlDm/sPmUou5iiUWJnJpf3EKDHMBXq3SaKYzzo0+nYNN6/UWf8e
jVj24GlHXbM9G8JcLV2MBlysjFd9pVNYlx+AlGUjMnnBxbZx4MFUnLVwp90/K7BH
4gEYeSU33d6m/5g4HzJED8uvnB+wWuSDUUx8hq6NG1dfAvS4s0+cWZmSiB+3gntJ
5FsjULNE7S3tQh91sfRXYTrEvLblM0JGgAZDK1yAwP/4f0zh5qmjQqyCAdwXAX9R
3zJie6uKmwUZnNNxgu92krGWeuJU1y4tuHeL9O3fzI/SQVRly+MUSRZG/Fnbdlan
sbWkA++U6EBOr13GhLe/W7ttO1v+o9/N060AhYuuFWvQCqthJMduZVmxAdZEDjUF
SUZAolCuokxjKAIbdbh2mTOzbSlbJHK0mAP7aeM+gvGPmK8oI7cXNXvigJyMQb+Z
XDIJi+LmX3DIAwAD2usKIe0X5p7JII8Ee61iEVuHVsfrZq8vSKWdnAwMT8xxnExC
5+TzJ4PTp1LmSry7MZmE7cPjm8kMvj5pLB1rwMywj8lhyYNXVioojIcMLyH6XFAz
0QAA9pLPZA1MzWfYOUBenbvtkwNQscnvUO8UiaqwLanYlRQSHjhV54jO2HH2Danc
wQsei5psp0BBugETxOK+Y+hovFfsqkSdiNyZ/tJxHqp6iuTfGJz6vr2IJxo2RkJF
WyeZel9fevA9CoBdd1CplZClgcrc0EnNRSguSxjUUGzMuPEWRUYFgbF6vnMbW6oL
AC/VZ3o01wMHm9k2SkFApSOgxx7F+YbGjucAjDGwNhWJkjRIonP9spC8vv95CtTv
h/NAMrGxS3qFQj0WsvifmdotEbSt+DetflyBjkfmg2JXxs6wYJvjBAgKZfM14TNO
Y3buKn+hm+AVUr89/dUsXfvqqLoUd/Y57NS32Ys9xK7dngQMbU4ZpOTlq135FgYc
3JJlumFU92wkgUQ85O4sF8aB8vE/IHBRV+imeAXyyICguJAsWyjAeDBHlk0w6M3g
5xz407nkGi/ynFkyQQWiGSFzfsHgq9TVWRCMd6DvPIdhhCkHyjl/YhhD2vMIw0G4
j1hmX0xOMG4tb7N1c1YDO5A/mZ2utq/G0yJl75iT9KEpSxAYTlrJIjg7gyte5Q3R
7ww8aA1PsAKAGXRrfnXnkBPc81F/9yHGD20rOqDgToL90UBv6+iMv8nX4ueMSzgZ
OrIIwxBSTrhtFNuEB9c0N9qsc4OfjUP1L0S1+EIiMbGekbpjt+/Bor+3RD0N3JE0
uqSdG4x+xE1oPIgv+A06S4IkP+3ZS50LgY4puvO9kJGJC4IXscjmRfCuAbondj0s
gPDbE8hYjW1aHYx6lqCp4ElgIQv9fHxVlpS/d87PbLn8drUZE293kSKn2wxsGNmJ
cUCSTi5L/UaQrXerWW4JUzYf1z3MVVKwLWHQa4pA1SlcM6F3e19pOvRe91gUIDnY
uI9vKsPsfEvHxiCj0GdKrRPg7nk2WHRIkZ1bluG8nr1mOBXrD/M51PcZqbxlAKRB
mB+euFZE5mEGtPmm/H3oJiYpbDgnlDhj0gVEbIvZ5Hu0Uoqh1efz5uctlg1fiJxs
nFWYpj/zGMqFGTXKDZBdzxU++fur9Ajprc73qsIKlMPO23MDQfPrcz/ijMwCFhPE
kbzPzt7dR2Z8voAOFh9/uNAewP05gPUS5KI6T8beIUYm/Dmc6nK8i2RAnGIwR3m/
N9lfo5q4RoMiZ+2tDI8WKp7zOS02SU6iYFPxR+RXCYwmzsRuZFhGtJgWVW9EBXsI
b+wkFADx58uWpgpsqBewbhOtwZcAJsp5zz3AV0Mcar/aKac3eyJMr0mHLdMRvT4P
/t6OQOUOueu+X4E6gjglZiJpme0FT6WtoYgU+b0uHWoDf0pYtJijxh8/PQuiV5ln
mi0PJG+KWVNo1hb/VtXBFA==
`protect END_PROTECTED
