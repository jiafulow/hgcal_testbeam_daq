`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHO87rg9ccwqozq1gSPGltDclw8k0z1lfnCtOwQh2+T1wNm720dE3E0etQ/Hre9q
vLjoBJ9jfAXeTUn9UfId/r8f6T38M7VJnl1sUHgBeLYX3CVaqGXfNxUPwtrIWuor
NyFNYGfGYIuUJ4xRpBM1isZlm2r0ZmGtzrLxl619EB21yhqBBtYn78U/pHUivCPH
AEhq/udY+4Zl8iRxqc4LjfpfEBEhjvkeOEzPcff7GH2lOYMex4KItPY7QApPmK3c
9DWLRyGikfeJ2Yr2Hv4wwKUr8ofQ7oHbujiVNOwZnNBk70QNWjrLNf98GmlAz684
NyBPwyi4JxtKW7rZNod0c/BARTaZIfNTEfqEgY4ZCO2KQevhdhss2Cfy9CgcJr2j
sxafJGTmynTauQqhqWa5V35P8JlmpfIDukmHbeguWkSbcFqOourpwYmF2QhBXuCB
/UVLRLOL0D61w4hTV0Ae0WgstiWjTD3Sa6ayGaaCQYq3uqFeGxd6ne9rKH8FV1he
u37N9za248/Geb8hqeLF4CJWOebLVuf50D+MqIUpCnKbhf78WvKp3uwUKy250SKD
5A/TnuatzW+xq2cduGFiKDZNH6JiS+YEWcDHx3W9UhENAZQCuZ/e7tdCFV+Dcqi4
8asz9mx0P9FwbJGmxuM1ESiVFtf+e+eQt6ZXmFo2lh3g5qaScanNrDtxXUAmLmyV
81TZjNHXivCm4lnWi4UyPqbDkCSfBI8692HK6HfYCno=
`protect END_PROTECTED
