`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8Q4IUnwMzMb4L7wf4Iai4bTrSX2BnYwR6rX0LnLnOnL8b+fx3IttKtTPTLuQWM9
4t7R9aaPaIQ7mR3yPRUNKOFTBNd0FKzlVFxkqYPAKm2D88cyL52TPweL4vVgyVUD
1pSGx2PDo4eYdnenY5pifb9VriD75oot+C/iFRIY2pYJvaTwa85DHiOS2ltku8Fl
/DJ8Lo0kBVP4eukFyxfyt6JxGcOmlkNOwjOU5Sn9LO+zHUVAP77RA3+3l6OrLQzt
3j/dD+c5Bwju/D8bR3+gaBk2O4UO19zKuemwXLnKNI6l8belnpx4xCQMuwV+uBuO
7Wwo3p4+gE4sLxrzEMY2+DBiEVjnea73jnVzItDvygBGj0yfSfhjA6FWJMOJ6qBw
jrA/XoCIAiB+BX9gQWrH+QVw+fO0CWinVbO+c9XsQ3LtLcXxNWMyCZe8fa01BdNO
6h9B+WT7c6VWhX2hX22TIKd02XD7bSycAg7fc+8xQJ4=
`protect END_PROTECTED
