`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
teMak9EvT0scoa7HjwDgTZwlyeUW66uZJDuE4qAqyqdwEvBRkmyZWFv5z/1iCgv+
rLaZCujF04FEWjtP5v0pH3JGQfkAqWrjEJSk++u2PdkwCM2frFahTwnulivd/WNo
tbseTIL1hQn50vbFAqR7oOLcmmTmTn/CbqeXrMgMLmJGSUSLbKpAAYWhwDzFp1ff
aydtD4rrAOMKjdculvUItcibTZLcROKBLo+33nDDtIv5b+oW42GUCw9TH1eMLc34
QGUXtl3+Z2ID+YegjPLtUO9h1OmDvS+9FiBbui8/KulWq3AAIFVyjFkO3dD8qCZj
BgGs4WMgOIWDzqnxfKbTfP0iSgR3lGpg6n1IaC6Z/ItU1MYaPbcGMvSLWmfRcOoH
pwGFuIX+IfN2yz/eoZgFk7ME9+Mc70I8p1h36vbRKQb1SU0px1uRzqIY5HFgOd/c
Ybm3GjUGtQtUZ0Ubk9UgEfcmAj8qDNkN/acG0VKr9dDW614C9zyIcKl5ShdcLH2T
926JDEoPwKwGa69KBKAngUYLk1ttOb0zk0U1IqOJy0bpNNnJ6QVCk3IhR8vJa21k
++ldPHXvNj/FY26/8294Z+pyQdZjc10VUMRbhOLeAMQ+Z3X9BMbli5ZaLOv/Ehr+
l1LACjAavznjyYVzbb12kQli+4mmWNzhCgt4LzW3Mf7oDM8/c/uvbuI5rKDrMFnm
4++67veu6q5S8Wp3a84h9/+Hf5ewGN33P2wDvM/oIolQH4gHu7LCPBMkDN6WXVjM
Zj2d4RsQvT5XKqU3KZaloCio6KZGsnJYKJrIomxbLX2B9UPfTEVfF8oW1t0Z6aWf
b3BIpXo0be+/fGU5n/srw1T6NtNj/McXVFSEIVq2NzQggnefdMvgzHHInPuRIorC
/L2M1Jr9hhCIQOuDAnOwElpyIUE2NfZiJPVHapxcyZMAXxfhnumXMHOvjpj+17lu
siUSoMhNwF2TE6ivtQn+A1FEApC5bNnkIN08a0xbtY5nK+WigDE02J+xAixB4I5g
/HRLCpmFmrwGfQcgprI4MW3EhlETI/ZhvvbYFdp68gA=
`protect END_PROTECTED
