`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pEXRU/6fTzp+nHBkJf43D3ZuQGl15r/X7vdJ3bzHmSr0+9Ra9huwmSnMVfKX+YpS
5NvdMN/OrnAT85sZ4Slc+0gUfanPh75PWkVDRkaBcq5d22x4bs10M3xxhpS5dUk6
Fz6n9I80ypPe3gkyVZcFt1Q8ZQpGQGKsWzVCegKJd1tIvZxsCnJcLbpdufkCsXBX
Q1CwSkTEG1pmEyPGAwtVqRUCno3QEZ+Sk0elEybi5hAqyQskpQw3bCOF+aHUMY/m
a7GXabtbR5O18PIHSBsm9ynCLkf7dscPYB2huHRXxYD41ohorvOAN8P94CwZ/8mf
6drQG6GM6kn7JyXFGGC9uZPsRHi/wrUF+txurfyL08c48Eq+fHaFmyRqrE/MrtMl
dsfBDPjJhxoWGrerK5CT3A==
`protect END_PROTECTED
