`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFrREwAuKV0uNgoiRJIAhWTNscpa82j8NVecmdzAsvW1ALqSo3XSHR7Nsm5WGOra
7WuE+8mfgOQJWinnZvkaW3r31J++DfeGEAlT/lOzMUklWjyrtTGH8lVVEjLYEoru
+jlCDmidX2XYPtj6uWpLeJQpR7nPJEzNjqZ/zX2e+JkzrApS/o9qDvG1t65E3yT9
rS8HSyNKwWZDqj3Mx6ZRM1uTpyC+yshRfYHDWaTxwszVvB+T/vOmjhAn9baYUHLR
nnmYxSCFuSt+6WS7xIFC8AAOd/wdMn8qpLTrXd6VOl+yzeAEdngtktrwSIXVHMvP
1uMju3hkGDC9+ZkGR38DUTiPV3pqPmLVqoXYt5rhrhtqmGBSBBA+2VEWK+thaayo
vuA7Pf9YB7Dy9I5V17k8miHEYadds1iqjMyeiHpaCfezgBki9uH1Aotb/3Mzh22c
yDK7XcOLu4F9A5QHgAGtgp4p8Qne448Kfc3/TNYxMXSpn4xbuzOzfLaqGAI1kWyj
voKVnYk7wWZQzV8MWufDrHiInOUFIL8WWACdwiHSWdf2UXt3ZnQBgyloYH21d2O5
9aklV4M7iyGAFPVC9Oflo8C4j6HLDvJjc9JCQTQlRCeyFeVmySMT29JE7JG+AL7f
++n2kq2ibDOL+wTXkLn/42n3GzeWqP/+7CImsrG9nXK/gxaSmxlgbjjlyGVpH9I+
F/o+PbZ+b+AgzwndUvmb9cv0n8GupTYIteF3ou5pS/pJOiIZJhL4wCvJCWi+NfMd
rgAp1pgKVQjDrhJfbYPn0VBXXiFfOSME3NBSqtEYxCNxDgAnYRS3gFdqiD+gej74
3ubcf/+BN8rvSunhVo0LJ05XFYqt4prCvlDCA06aMNZ6ybTlWMfBCCna9GJ1tMB2
MdW6Pvm3ctfHHNRZaSZDUGlelhmZcqBA2LxLWyG4eM5OfAZ388lZQkkTvXj2q//c
FtJq3coqU4kZHTsgqftpIqINAKNt0JQwBsuoyV4vDjQWtwa/6+VGT8HSfnAgBPeO
qYf/83PCCb+IrzvgkkM8nlkDmabXz9X4N8v4tcvRH1tR2H0PKnY+99KynPZ0bYEQ
oNbTThsW9nGxPnOTpbSbvDnqpwZ9h92GFNp+V8Kp9TvIs+3OvX5WkPheooe7fGNp
kfHKbe2GPodebKN4TB7iqtkcvh2+AuBejiG8E6ABNMnXAo3PdWygVbRV7h3r5Oqo
lYru5XWM4uxogDe3w0DaX+Eqhbbf9NQgEfsUmbKhzHuSuiJuHRyUtOngSaKghkMT
CGHrtD6qw0PUEbNrhyQu5fmir3wgbjbQYkvSJPDvraYBw6PvS/lXGRNfP3j0qUf3
9EzcPRp8ozc06DrnVcZEQ8V3mIydPoMjFjGinU3edHp8m1NUN7rMrb9AeINqqOcv
/qkmVXx4KTJsClrT3cBJO3MqlQjBFMMIFLcW2N5D0Kz5F9InIprrbGkT6l/MY/AE
gsjRChRZh2oF6rk/HAJdTvcFzAXhO5lZnbaSHz1gdtzVhuT6XigkZMx3M+3RkJ8l
3v3VRRI+IG/isVMIHCV+BNLXulVG0B8mJ+I3lyT4mxkSZ3iPf6JnoHGQRpO1j/jD
I47vET4WyNNnWUuKjLiT1R4dWbQPBhZD+3RPT8VQiPmgbGhafe22rAnjw8ST0NX5
cksrqzhX8rKCnK6ZJdw0HxZKQ1EcAWnksPpZy5T2my/a+bV8jHrRTyIQhkVkQG63
hMTIqrfB5wLp87UF4OfqrRbRjgRugcX2MT9gjM8UcWRP9MJDlhKH1ttShvdBKSAz
M9jgxLgzFC3yC3lc3K4p6LnXDGtl/SF948UmqC+3KJ8xSrZaPjgKnS7SKnr9GvCb
2jfS/EUEel7434ZO1t7F3tceoeWv9WOpDwKYY2A9WIPZ6qr9L4hbyB7N0T4udYPm
53mv3JbHL82hdMQeaQSysfM2MAd07t0pHe0WLwONqW1YC0MxJTHouWzHMkrmDJoo
HyyigqWmlKl19ZK0VUEkvNZf31KzSxVnl5BATnYZiyaBTSYcqmlb0tZTjpP01Nlu
JG5k5kpQBVvQYrNd4hZHJU0FJP6gjMtd/esStja6MV3P5oZp6q0nlryv+2t3KepW
Fdx4q89Hywndp6Epio3RpBz/EqM0X56fT+4ORIeF0sF6CjbZh0umvM9+I2ZZ+Jsp
o8mEwyHdOb+dY2AzDJcvR2xVkuyRJCYDvKgVrywGXHM0Swgf/Ed1VpOB1veEmcYq
7F2sdS+zQc0PaiYulX9h46CBmHDhXTYLtA7/GgLDAtrR5KK3FGUnwGYwwFz6aai3
rysADtifKV9GDLj3JUIQNEvl90UdW36UpX97uC/PJRkzo+7jWW57oIvEpBakWYgl
OF9LsvvD8BEh/OZCq3pSDuyv7oIg19jXOKC/JT+zAjkVw8geSOrDjwVVoFdtSHhL
Jcc2pd1dtgLV+N71TNiPHktF/STzlo6qGtLTYlPO7Lusk1ZM/elxhhvQZOrCNQZI
HhWNZQrOT3Z6b3e2kqnwjWnDOaO/QOAs4d2xOg9MfkqQ44v2qFglh2rrtfaOsvqr
OuZxEC2M5ZpYu0BvaiGAGXNVbjAOwPCkxENSXQ5j0gMk1/pRZ1cZtN6Mms9UNRxf
jCcGxMLBG/TYwklPwlfM0cqM2ZBoBBCcF23mfNOEPrFVx/aHROW/Yg41Uh0Ynek/
9LgY11Wn0buc3drRGMkDSpgGPS4oFVeO0+OhSVMtIy8WGFIyNEoD+8mDq/rMSNcr
0jacQ5kIG6/bSZAEQc9Go90SVrSTbl5xhboH0MbVuZCnyfXmRLx9n+DTyK4W5pJm
ocK0oGktXbsVQzwCweWM54+wCLqL0QxHHWbHGJ3suHnHIqOWnurGq4ffQ5wA26mA
FC/1NJdRMYhqn4td1F8xlEx8nmIpB4llu0zebS1wviW4DFkDw7ghwKF4RNASLQ+b
1kuzWpMIWpZNKeY0oLWyAtnZgvOhaKpA1LX61+1caY/VHjmEqGGTj07dzS2vY5wx
NJNSajkstoVgNimpIyB6Uba191Q1ssT33i24hkPj4nvnU/DNb/2qCwB47/dk3PAu
qY24vIElAoo+vTDxDyXMOSnMSHis5Z4eTtn8RSMhEoWeZ6NudagX6bObxEYtbq10
Y9knUX17i+yCbfhRZSRk4h0PbjEFP9kcSypz3kqTqzTE7NmvddydRQzAGPetec3J
czN63Rj242MlUxASDkI2mpCxHtfmccfkb6jR9i20f7ysVM6RQeyhW7LlPCsNt6BY
7+BDrFoYsq8k04TF2t9Fq3/AhljzS+H9LYQmqtaGsjBVAbrbHk89dRo2LFt0yGfE
I5ICc9DEAI8rhwsCBajX8N8p4qB3A0A4bFG1oy/WCZjhO53oIo5MYHmxGgGFtdLG
7sa7i58PXfUh/EjQ66pofJyM8nUOeFpkIbPKen3RUcD8eShM93hOUy3ns5ZQw6g9
Hap+Ggc8feh6rvuSMT4W7b4MgY8pkFOJ9aQMZq67EgaA4M2WM/cmX+PxcYN51kdY
ByfWTM1PxfU15BuUz2tOIxrHEg7wPgz5f7Y6/ZAUnKCvO/WOqXdm4s+A+pEDT2n5
qEn8WSQVSULBic2AmlekR47skfTF5GdqFyHAnQcU7ZlI0dBj3T6mE3sdUtSJkZCy
c1q+cR7N7TUmcE3H+QTocUFHdr3FpQFq0LbQhDK9LLh6b7vqlix45GQCPdO79igV
czoWoF6tXLft5J5b7pd3fBcTBvGKw0K+WUhsUwWrSXe95kEw8HT78vTUlBkkDu2d
9+KCAaGm3LtjSnV3xS1Nh7GGEHAJqPd9nk4ULfoVrH0TMZdQ5tV8T7Wpw6wFjoUk
RjOTFCbWbSVhvOm3nV1y5gNUWUzAOc+o/94AwNyRJxRrxWqbJOYO2scVGLsXSBKn
+OrAsAOTU6sDyuNfJiHeGFcqmPeD8xU6dtOl/nHTc3P74tvq7jeraSa+fskgvQpf
0KEpzl7BDSTBgWk/76g9meeyOSXW2WCN2TivaBbVxudo6ZbzBsNJTHX8UU8Af3vK
7ZJRgyjh+xOHk14INbqDQ0lcKWpZnOmABgSD0wCQlNPES1freJKWS2RASnb3C8p4
iwiaj/ufTr9D0tfcRG8eTH2F84sPCBem0YUtEdCZzKxOwC59HCv18QPoL/wUAsiv
sXxQUpgg3EHlhlxKpzoGvWY6ffwL1U6lJYSr7Rt4nCCLIxN2VXsPnMQ6CtIJdSqX
LjUX4Q1bDg0Aq1iIjtEGCD46fGXRkpu9jGF9tHlxrMVS0gL5aqqEwEGo2u3yoWud
ADjzWwsUkkWDF3mj1f0wLa6ZUq4aprOgAZ1oSaNe/iqR0ildf/9GAuCheYW3HUBh
x1616I9n1l3AGu1MMToSS/bq2YXWg4QTGkz+y+dEq2Iy5pclOc/GUDwFuae3SqYg
ivu+PAi66lnlpcI9WS4ujEcEgYFwjslL9a/L1wobSbk4mcOSGLyZHxMoRrCl3JgX
unkNjdVqSe4gL5CxKW42Ly7LRbgyWIyE504D2u59HIOwAd+6d/1sTzBxLt2xtulr
FUkV9ya6tngxR5Ak9pyx3VnK/FSX/eh6buFTzlERInDExbf64DhAtOBWuncGSFkJ
J0+udWV2XLGp4jZotarLzLrWs/vUYUNgbED8ycMQF30GPlZxbl5sJrdgsLV0dPeH
ao3TnSZQpFuUjA4lWkPjuHSDVF3IeCbwfk40fivPkXWg/WLScspKy2AepaaSt8vP
XqbGCB+vEZbn3zkSaWNHwslUfR/oyz8PpXmkwBnlszdL+Htrtp5l6/m2eNHOD/lk
IGjS2CiIkeQeF0eya1ItPdvN9h7s+nMFp3hXrM4ShbE7M+R87X+kyCaN405n2cjz
AUkInO7sfLQO7wQn1W/lAsuQn15vrRUbssHXOFLi4msoYfrQqcCqXMzIqN3uoX4Q
ZDwA8J1fkPhRijCmHRoe9lvD+hMS33HbBO6h5fjC6DCLPy7xSu9bmOf3F8GGokLO
6gm9vIOpo+K/m7KtH4JPisG5pivI3jFO/zkhLCS8YhZ1V/rvZT1Dh3HjeFDJhCNo
wPM1lyBKaMQuclp8UVJ46j2z4duT1E4YNhQs+OPSblPBwOg3a9SMrgEOeE2d1xTm
V8Wf514l7iOcpXEEltEQjPg0q6Y4PzwQj3N9/rIqqqd6VnXEY8mO3+NzlgbmwNjh
1Sy2r8ORvnwax54o1K4qsChIVF3X3eFI9Sk7ZvV98xqaNd7BWM6wv8ISsT3Te/pl
M1ntgvYM46ExVruaZ3ZyCowewl6+DAVogFy/FtvMRw4cX7iQ1rbj3vhoOInySD8q
5kP02Fja64UIRKmUFuCLu4rAZNpXurR58jQ3WkF5XALt5P/CHnexIk5zhatVp4+/
aUUcKglKCkfG7rC1FXyJWvT5Pgv1w4Q2h8BzUkXuLOCFoTqrf5IBVL5RbMXqttiT
8OApoYikLrLNi5j9nWXEiEUZ1RsnhKtGn5lLkqWN3KqVMxI30SYuXYl+98hfKktS
iKx3RdNYCcL0EJ8dEatUhH6zTA0XU6y7pI9eWewEAajpcACyU4//W0BNNG0pzMgH
DYIxLhEM2URVovtX51bgPEOf2qkj8TW9uo4KoAYG3a0ir7KjrL7VdEH7jm+Xtj6n
rVzK/w71MPqUNwJhVfURx5E3qB2nvtttYfbp2ZO/6bmCHHtUARr2hWfIa0ZgBh7I
V0trQGJbc4/yRJ9nMLeoohN1zVdwMPhvYNQbI0aJL8SZU9Zv6WAI4dA6Sf45cAuK
IbA5YJejszGEHCwaeMsX1HD2na5A/BBbo+Am6E7xARrhMGoMoyMrnONWTY69mnE9
aQHIQd/vIU1magbDpSfBkZXpg37Hcisz3ksmtQjBZeinwg8Oe+fHxGTrSt3m5O9v
p/G8t+iR7aNJnERWUG9Zjr3MPzALa028Jlcu+bQwNAw2G4PNRdS5fZ8kCJBs0k6q
SYPiRuZUB4Q6RmwALdFiKpdFhVrPCbvX+6dTpGJOPofu8dC/i8n+Lyiy3WJTGHZf
gXajWf5mN18UtmUOf2nPx9+gK5sni/sbfZzXmPcmB45RGyvAkaq2FdvtarmfgQ5+
WuzqBg33I/hh/qKlHSXFmL0A0XmxaF67EJLMho5jBY/jjtUfXIJxIjhlHqGvhLP2
aKuOtqbQzV1O8O5gAxelRrPirOrulHugbAcs+oarQ8AglZlG6z328lLVTBkJxj8f
FArfEAynSDTBpQLZm7kKLvJYKdzr7OF/kvO6qX7f0PXaG52FwrqTz65JryD6DpE6
REphyTJo0m4W41ofdEimfplhlWWDUkGAjHu7oTVXdTyDq0CVsISaicJlejStxijV
ztmCwir9qf3kt1A5h83z2JtDrEKQcf3XH7sHmrjyxaZ3WYyN69ZTJVeu+FHlyU9Z
G0sPuUkmhMs38q7ErnO0lNBVtyFVICeB52qMwO2HOd1wwXQNqKX39AnBJ0lLmEyy
NqsKpZ3cspoTTzmCxHq7s8gNG+fPmd20gwVFm6AXfV8Nzz/Kw5c1kJrdI4f0xQft
2fp8AelCeb8pm7nKj8JJYwHixrW+arSaUmtAJqORVw7mXRhsKEP+q9x5+WIM5bNs
4KCAb7z0Hma1kv42h9cEdeVX9WgeD4LomxWPxQqYv9Da7hfWtaWN0e9pWr7BkjMc
NUbZ9SFxqdClGEeB6GGP/gVePVkyg/sKEFR+FpstgvUB/Ll9mgBLLZw8WxaNkPAT
mrg2R/KYh0r65Hc2WNcqLUeHYQgjbIuVQKjTE9iAPZV/VHqC4SmV9LsrHZxUovWE
i/8TdTs1EK2LMC3kMRQLPUBQPG43SBP0ZQMc0bb8FhJ2O2sks73cy9hBL1sXr2/t
1HV65GA03akG9PnhqxAzBTK1mfO5LF90kfLR/wZFOpPQdHFMIBpi+19r3kETAZZY
9NpezL4efpaLsRmANeGTcRfF/7R8kFnbRz58yyHfwmMXSCFtbSqYx5lAvGnV3K5l
fzoOBq5DVfGKL/RTVQ6BkPzgaA4v605nauC4r+hoAP4ZIkuBy7pzgJ/+utNIz74x
yH9RLZQmMZ20WhiuG8JzCMs32ClpkmEUVErcsuY3+lxQDG18hCRcUNPgNiuj8COf
xBKsu4+3H10kZLYSxq2DwqVbBTysoi4mGgxhvfQKVHdmZS6DUKRFWzc/i7lg7jHc
3I2Hyfp/AnzQN9h+Lo5MqGeY6hCDTWYNkWVOshWLx8cJh50NHNq2PWHIEcZFltl6
WmXwz1sW0Otg/ibuj5Ufvz71ZdpQbZwhpxb0oiNrn8TeQHGYkSaAu5exNPI5kwnR
b9gIQhFToFbr2TZ0yBq6s9eDdqukLjte4+m57OGuis6thQpsXpwaMmV+a0AvKoxk
Ur7ojMoSk4dYJnohAz638DkulCTl48B0h+G4v+WG4o8oL4ve2CtZcKcagzfGoxq/
QZOcrwHU9+SicUYt5zFCspY5IJ2QCy2ZqMlvvWNkwX/3C/1eT9LCVXGz42nZNEGo
Vyk8Ng+2+A25mLB38UiuTl1VptJ5akKzQfNC1o5+iOOJPwzVdqtcr4PA6C7w/byE
pfCXVbfMkXp5fvAMMTaVRzA2cjMt5Rc4E7An64L4dNLCM1glJioY2r0NJ1EuaQWa
PWfjSNB5ikTf90whvWzSdspDbepw6y1vd3ITueAOXFvPYVUqC+GhKwr3eK6vHWgT
1TO7pUDwdFw+T3TK8z7QbpgkVZUU6JaVlG7C9lapuxZqi8nffqUt3oPmS9lZiZP4
NwvisaRU0cL801Ff/XNyarnsMImDBu/AdeRuqM+hoF/NRv5IHmhGr2ivydl3kk6t
ZXBr8Hmkl6rcIPu/Qm9Q+iwQJ7M4mUslkKawcdu5IkWhFnmB28Ag8t6w7ZMO905n
`protect END_PROTECTED
