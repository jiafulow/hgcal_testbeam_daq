`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZLq9Wwn8Mi0qZhwxEskuUcexwd35EzNL/rbzGs3xmo+7rmz+9AnWfM/t+SIUbbQ
G4GSpYzIJBpIDs1JjO+ovbtc9LAZZ7gRFcDM7uz/hkdH8KFV1mj+MDiq5hCSuJiZ
n3T2+x2ePJJTlMHWjrcGKUg9laCSc0CbRlpzruNUvyAjfliXfMEfEzkwNTiyiPoT
f95nnG38xBkxt6Rli3JxEmma7mJVbtgE7BJ5s+o3PgSPXAG3uIgNNweZuo2fdOKr
33lSodNJ32Qg9+7BFyVEcX7qHb4Qj4wHf99IFETBCyUSiAYTMxI9bfmSqLvIFo2t
HdH7Lj1G/hVeLIwOkl5qyhAXCAiTHWPEihGD5tg8Kyrln4CDpFgDVae0V2l5qK6U
uUzZotnXQ30NnIs3rlPxU5eYwwpn6VWTpxZ3C0Kwp97+1sE6cVMlaHCK9BOmpgkU
JxXnRg01z+zFjWdZcKJZPErSg5148MYeOXCu0j03j2J1LWvi5NqWRh2qjvON8Fdf
nYMA32yZtOoD+/eYByxfLLkpjqTiUCAMzeYdD1xKKakQ9dX69FP8EhjBC6hHh9hH
EwYW5/o59L5WEpgiNNVTPF8XLFNR4zRJ0qC5WteKSoTSC3dKB/ovBE58AYrbtJhm
YegNv5FuazYAu8AEPox9vrtSulRQLapDHmpTp1ATSYGDSTl+8PqZelJGzx/PHOct
9RQWB29ctWXPaj586ESyJClyvVosYOsq6xq4v41QnSN8sMIc3X19O2W39pMsjur1
tk5vfLkyhpHUGQwzWynFzCJA+Yu6kiHz6bm8XFW8wq2qlCCAD0xggEdSUVaTdkfC
NJTUi3ZGQg/qh935at3oWNLctJ2h4EV6Z3us0me1Rp5X7if2Jotrf8GcPiSwsnwd
eoOB7vG9GUWNoXYaBOOPQtzRQNuDwZBNv6rQnR3xGJa8iUPCeaS/m2kEiLGqfdtH
v3KPy56AumRPUP1MMrRxeJdbQ9+syjbtsfOJp30zH7Iiv1cnD7C14AExOR/nxCUC
2ROot0sGAUK5hKs13sihAi1CKfPzWhag1x6sg/TAtMCa0r3Bq9zafUnNSTc4Yor8
RB8aBXP97M1c66++/BnYZYbPdHMatLB0ZQxPmcHzdoDHtzVDTRQiRqSsbg3+JXsE
nBAiOzcYzEtSTJLwUd6Girr8PTRJ4GGYLPAa5jxNKow=
`protect END_PROTECTED
