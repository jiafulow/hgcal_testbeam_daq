`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iA0yoZfth1ItOjMfFt5iFK+1FNJlL/VW+ncVJrkgjURgHSjn90v9RpofgqxKO/oe
KB6q/oBZZhLE1SSmA1KvTLBB919pnVFMYmjud/MaH/TreW8JP5V/Ngrvm61/MFkg
3z5eVDojJojZ5+1xoHQu/+4hUEO+pwmNshE/SzS8zVqiWO8B6rYwttkB9OxTNpXo
C1BV4C0dMVcF2un728aNtLwI2AR7mtsKt4PCI+q039leLSI9ZXBJU0ZzKaTf9yLM
/bihx6Fn7g8IXo1PLZ8VdJYgq34pNc+xpnPExIcQF/TjFSuS5foB6kVrxBbTHC+8
P0RUMT8VqmMoMa04N4XqTseKee5u3bPjf61dY2ET2M7/pe48/5+BqTJfDkRCsFdy
+0dZTWQmwUC1sOXLuR+c7gd2kgof/UCSuOziarlo/PVeSUGxvJGzhou6K9kueLMh
brEub13VdN3saeLOxoowhwh+5Zg97yghsDr6DLMEATTnXipwYjcL5MEPywTkupds
b9FRiBTRWmGie9inMqxTlKy3INC4gj7wqfJpyN4yAeAfu3E3Zco8xIWNuMlg+se6
D8sfz+pL1rDOVolSJl2VSgoRIY4MgfdOm8Wr+2KALwuUIq4d+c/XEY07OVWJ96wp
F2o5dzTYbu/nhJ7FqzQP28fa6NnWbEFgwGRrAMKbWAepUSlaox9XSjsxwvYoHOgZ
sW/rtY90/8BfkyqyAMmfzo3NedoTWxsvKm0HDJ108m3E3GvGuIbD6zgRvV0Nfl+t
AGpmmJbE6WlEw7R/Ju3gZJVvYWS04ECImjNlHOpSiA7xy4sPy05caNhMSbZ5PON6
aTA/SZaEc2P7qSPnqaVV0zqUz4h2XwWpcKtb3obMfpTEJZfu3KnCSL60KOEDvNfy
nVC9vIdglyOD8CcD+XudgD4GXD9fXtATZMQZHizjf7UWiXSKVyqH1Blpx89PZFvB
AFYbXWzZsSpNHLrG+gvAELfQtj4uIF4pQ97QUBuR1HCVTV9kXx9bP1vC3a7Ituxf
Qx/IHcZYCY+JBQ+UVAXCgrQYVVPj9RNe4Pbtf0zrJRucXo/GeuW5hZI08XuUUkrr
7roTPIvi9RmIZahxzvfpTLzJSl9ZATGOWheN0VUL4qBaACyl2pUe1dIgnwHy0DrI
qE+7glDIIW+y6EKcbyQnz9QzyMfeWy1rNy5iCaFZR5mijE4W+6O67K7Sjq5R71iD
uHSiH0YdNJ4XbHSADKP0X4LKfYqMY7IE3TpHZ2q8R2fNcLBHwbXBhcVha6MvExAL
gXp8K35tCikQzt/4SsXwwF3npjvIUZ+WfsMYUVA62sIYgzPM+mV0894iX0av/Paq
u97891lUfW5L110tGRlhTqQuaDrYMWDojuMi+9/CN53BbvNxb3ZMnDQtIkIYqjmG
Bc+eIcyGhmKCr2RaeIvzbWXEn94qCOGKnu0wjFBJJv24Tf+SOr4TqjQxhH7w8ftw
nzSRDdP8xuKhEeYp8RMCaFDOGbPh3gCtz55G31AcgmAUsm+gXWdH1uhiA9UxUiJk
KJW3b3BWnz6zuMZccRP9+/7zBVFjq+W3EmRVYpWj1Lm2yGqhjuZfY9KDRrg6P04+
76cQocscOeM2vgQK8j49pxn8ADqmR9hzeIt16Ax0YJR93Fhj4aeBM/EpKPDviqJH
wct2G1b4aBnMaoprZsdOiC7mvEqACDbfIv9OpqeMUpiZMjwq5+YL8BUyaQUepPwl
8c/PRVO95csfxoWJhGDO3SW+TgF4pYXQSzrG8xlVB8EridCtPp4po5j23AAVvCel
3Tg70iszMJL7FGElZT2D0g40MSVxTq3Nb6ihkKrksHT3N0yNlYZUw1Yk8oj+4bo8
yBQWnjv+cIJH5vlsnEunMJuMFXTNcQZBjQyo7PdnVW+o4tD9D/M7boXME8QpCU99
dkHGnyHH0myTR9GWE0tKP4PT4CEkorSgJprXTBZstZ0=
`protect END_PROTECTED
