`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7iwaQqCvM3NG/oBn90EhFXbMwy4BOLc7bX6gNvzNvBP74gwKaoAdBLg1S1Skzbd
l0Cs4gdKEkuP/H6d5BknNiqMhxb4wXIDBXUAzLygAT4ZWNZ3sh3O7dSH5VWR4IYY
waR/OH/dP+u7WdWusHZV2/rRkbO8ozcJ6K75XStMUtE4E8Tw5ac1enjMsjJNACWq
dvw6OG5qbFfVwuoJUk7Iy2GzwsxSk2cB7Xb11BSyScNFABkuwypv2yq7IfQgeuz/
HUPckQKkVyxRhYU3HyVEyIkn/3U8F2KVg2qUvOh7RkaIWF3OyN73gcTc4KZBulNy
CFwg5rDGOi/3WmdeOfSGWfYHJFDLNuF41KWhsXOFIzYbP70aoq5t+fE18HM1hJrg
DZ2dbpCOiiUy89QQnpGa3H6470weYP9CJfegyT6VgK6YW/cD+R2ASYRU6gFOUTB2
oTSphOZ7ng8KmayCO/tHASwVMVIjL5+h8+rHWJ56GWd1WZ/wCKhyOhjYvMlqqYxh
tQs4Mqz60Py1DGynKFmrsT8itsDT1YGfRYZFi7HtyIZPEfamoSGhdoMqg96kHELM
I5bmfr4GZnqqtawumthmKQXkF4TxUaEv/NOji5ri0ea9u+Zj31hahK1H3uS8s9GF
u+Dn3aBRBMfOCCMaurNMMDQ4DQGxL4m0aAWW2TUaogFr0zyI80yHhNw7qQ/k1QzJ
w6PmArX9W/jWZPBgbdYSdR6MvOIvCtvojZvwZDEgcbmpwTC6qH+cia3hnO+ORfkE
sW3uhll8K6PB24wBbuSYJmVi9iiXta3LoSgUv9ZgVlDQEjQgwDKaDYOWv1jSEaIO
fAri+hpP2Bejy/dVPZAb7Fg7cOG2ppwTIG4msfPuZMR56YBUkwtV9aFvGb+v6LPw
pVVSJGjjrLfTuzV9oz7K9eDAFZRpomBX5fPkYQyDCIfSQhNjfhaZB/HNERBhmkJj
XzRG0WyZh4OFZTVJz44YFIdu+RmF0nylvEiD5VGDaHEp1c+6XK3K/IAytBCPOphR
9igEishEiWIAyq0TNT0pdaOSo/11n01jcNAbrsj4tomQhPFQpKLsqWgkKQSuCHUq
GeX7AzSOE4Rzl6ISyMS010TNUKHQ1y2rMeCJoegl16/iE8+Mc/DrPanguf6+whfn
o5+ZqHVLOVM54Opq4Xs1Rz3tbFyjS4uPhk29F1bGhIgkIFZ+C8siZsD1n8Tb3uRE
DvUl4mI9ZJO56Wb1yJp0lcc3dPGZYsBPvI6BmhFKKHrbTJaQ2+jQtwOoOCUhuQ8C
s28BQ8Zsu5NX80CCJEw9uPI7woaAfTq+MFSSousq9Bj9au76Gx9wUTRQWcPwiUTP
FAl6cGAlFLh89ypa2fBjX2trC1bUewX/HnZn4OaPt8Sk+4UPfSFTrBXgU5uR21b+
qH1iXSPr+xttRNPjzEehqWgl+xTti7mUtE9SnjU10/MCRNoRYdScE12xeC03p1y6
Hu+ZzlNP8gg7m7SYEPB+09/K9U8AQI/YxyDSpvl3tn5jlAiGzd1p4aGOiNdd/k/C
8nLFfO8PWSPjC3IvdYR3xIODh7NEgNTRsIieWmRLxziiyXoXYspUAli30/ntR0qx
fd1X+TrKBZGUua34Py5gC7Mh8kDQe3WHHoALUmo3Z4GoCnscEXjPytghmVIuaTky
XfTjEdSJhjewvQah36+u+aXy48b2PyiN+rwavwinx1iYgqCbHwmkceDtUdqF1405
bMrFStOUabckoQQubQWxhdGA8UUEV7tS7FgJ9fP0Fhp0zVz7fQbdIMWVnizy/496
BEcCWDqgiIF51RQIHJRQPOPZdODaQbAm/Zsxmg2TUC3qMzX+jCrnmrkpGDdImyrt
7saXbJNLHJpKg9IwkGPeYQ==
`protect END_PROTECTED
