`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+FKrwqX8zXuC1BVbkVB6oH3oAyI7OTAofENEbhhuAuo1nUzX9eRNyzScScOLugJZ
/ouv1VSh59NoQfY8x3aozVJlNx039JQxzDdY8owlQ+SEpaY/YmbfToJMZUAWhq3n
LWKkuCbKTSp12csp+OSBONWO82Enj0Jie+CkTRbYu8NjBEi+VTqNmYBica8oFEeP
wahJUX8zYOmsytRTHKPJGa6v9KJxmqEHmMpB1OA3z1nl09N4/+N0cCAQYr4IxpEa
kkNIY2NEA5WRTw4zqgN/QT/pkglJvmlRjtDO3XqbTFKPhSnZPaCb+ZNz+is/FJBf
gMfLScjCZPY/LzhNZWZzCCDGt9MZDwmUHKOVqJkDrZ/CeO7Y2Y5HTeqZdMfhPlwE
ETdrlYjgN0BbWX7jIOoQeO76HEBLiJmqXfEV1aNTkhf0cVB59Yi9n2aeDqE9/S5d
L0NM/1NhYu5GswHKfde+S6avowUY2VGtkE3i+blyzcr1XqlDtbRcmTLKs+Uy+Oqw
zitg/0hxIQSzJN0c/CH1AwHSyJrdk//fpPYh6DDdVR5azidSKDsDPWyfuPhhpszK
uzigPghtYWEuo0jywUEExS32e7q/pYtYZQqPk8I4g3eQwAbx31rq5d7VgK/qFgIi
KpDPwUWXiI2qF/SRCfEutKb+eSxE73dugS4kt3Lq4BUrmk5ZR6zhE2ojZ4Z20vAA
Fj81unn9tOkWReEo3NyOGeFegem+zYiEeZPJmOk6R5EOVZQgXCLk1Rb8vWXgJ5lj
mIG0YebzLBeSquC416aATV4nagFJTDvhGvdzAKRhJTUpqRI55LHeZgUqBu/WVfJ9
/atzKIc5MiSE6gnjG6QVZOQaYWIwAPBRDHMXQ712vN+t6FjqeOPCOsyycV6VkJ5y
I20pwzStq9QgmZSiPfkm8fNCOfq6Dz0jxS7mtonQ46L6lJmwl9OssbDP2ycCL7T5
dU9JhwpF5ZcCDcOnvsTDtSTtR7J6+7cc2zAUY+WtxjXXqH2qop5fnlNpdmqtSHsc
3iS5N6ShRi5GlCzR8AEE+i/G8BhLEgYUiVwpIbbku761+cSzPvLF0c3ysE3P7sJn
Cf6dO7KZOj4qvNSs+g8/zQ==
`protect END_PROTECTED
