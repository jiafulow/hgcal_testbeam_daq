`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gwoo+s6Q9qpGhOYytqN8REZ4OadgVADH3cszQIiLWTJRnK3CCfx1s9pUc+6R0Pp8
AIdimD4mn5RWtnXSnsn9bV1aF9Z47XzV7m6WiVYkEgy3Wbtxm1Y8IARHGnZSZnmk
fQ8PF6B7+Kr1uhNFTOeVNg965A7qlZhG71RWVfJJKs5SMPJvkSPiirIIZ1BJPtxJ
X1hFY7+ELrw3LDbf9ab+zX7+z0YR98V9RXJ2jcwJ3CQSF2YlUZDydiGYgfT9duMM
/NIkKdibh7mVGrKJp5xiT54MhbnqJVm+0qQw3aDbSK38l4oqWh/F+A/5OJe8Qy8b
wVGA0qEf1ETtQXkSThD9KCu9UJ2H5vbV7Gzimo1vq7yLSBWw07FWODuyZdxYUY9p
0yik14bhOiJFndh9IHfSOlnKd6dnaV+g191j9THd2qV4QNQTGGv/MiJzPLCI/V1z
liNJeX5UWbQvWytDKZ9mqle92vnaj0Yiz/LITZBA8DuVCIRyH/aOIErWfnuSQ1uH
aVuN2zmFeECNQcImYiJ4v/86/KdLFavmiuAQkjUr7fWBsdq9gW1DR9BeLN/iE2f7
B9iugLrg/P1YdhRUXuYBM/56XM5HRwUrt/MFQWIkJ4NhSQxAabMvXrPM6uYZHU9r
wu0eDU/PbRZDyUY4+IYcmm+Dx03kbqnnunK+BovB1HOPiHY75k2ZPCH8VfP7yhdh
Bz8ZGjegNGtI+t4C/PHntvNPIFhQcEzNEe+bY+OGzl57ho4u+ihCbkQz08ix4on7
/C5l7TOqVfG5Z5cBiuHzRBZuxo/KDMGR6CFO6iudbuyzppZldTvRoKxcXm/MHuaj
b9ju6j8yhieqDzBo27jGyZCB/e8FqpuwVxsh3mBVQO+PvTyIqYyvMFB57qqIsxZT
Z/KBoj5GcfAR9krxg+Gn265fkTafP2tbTf84v/ZwRbap+HDeMV6NLuxJ9jm6NlTO
8uxFUYrmpaTtEX3cjagjEuG4xWjTuQeR2K53c8kjiVHhJOp9ubIaSYHD2jCKSCpX
aaS3QBePriZChd+gVEdABfkaWv73UePNRLdeY0Q2hgCK7L1hu95QHLDlrLcsbXer
5uzhsJbvLsif0vSRxlskYGR1a+P/J0IpR5wugaVw4wtmBD500wABXCCBudXxBoNI
dJh2ELb1BHdHZS4yyez6wfkp1MEelvbHOKhSRDUwf3TTZty+BEziC4h5lQbZZGUe
aTLadhP1N1FAD26BOZqWsk9ohHUSKSJjRKwY5oisT+aygriPX+dMdaxg4CzOQ72G
1t4JN0ZcQR7lC3StGuWYwY4mJO14lYX/eUUxwGpcxsA+zRx+7qbfrpUFeZhZNsIS
4oL+Szjn/p+xYW8nPQ1kOlX88V6200bH8RhZZvqOihiDOd8yVgzG82/9QMHLkv2f
YO343yZz+wpsssCWueajyh8mzYBD5e6WaF0c2esF+lNKljCpOVw7FVcHu1N77BK8
+sNLetgHz3MLIKO+anbFzVXAsroBHUEsQJhsmawdCfDZO5XNTKnmNdNAY5KPBFBX
uN3NjY3oyG0PZmHM9zR+Ish9SfzG6JtUY01tL7SEcc5MSE66sM747WD2DkH/X05j
BqmnGSyLbeFF/E8e7+boDxHCIt24lo9RFhLJFJxmvGO1ifB5EKTwz1200LlbCxL9
6uQrhUlkcoKWQdsO9lSJ7d9azDHjaqiD1lx2vssG1sSiw2CkkddHHHrcYmknyziJ
yKTdvhCcQLPVAFRBEfjTU16ND7/jHkQBcwP0QIVteEJhdX13j5pX62yVoKGLmapf
8/WpwJaoAdI63yDfJpHWkN+Hbm5rglGsjH9oxBFWZRwEIVMwDZwN5faVanFJGxpH
Z0QMHLE+hl0VifO9DxY8ug==
`protect END_PROTECTED
