`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDusCYHee0S0Hcn5a0M7b1+74wnrIM7qJGRvxfO7EL5dfYKRO90xE/jJD6Nj5/Wf
6SSUodxy90+1GlRkv6gZayR3yBtoBy3bWFgdbTybCVUlGLoly/ipmFX9MLPY2X2C
L3LkmJcSwldzqtpGBcIL/o7bNZIyUR65UW8y2T5aAn8Nt+zb65uIZZ5dEj37Ug1J
FgUFmwJGpJulnvIQJMgNOPD8w9q0m14eSS3YEwW2GmM+inHauD3iivxhTgbMYNTv
37bMPBlVNPsD5vbK+IIr2ccZZyvDEhCQ8s6NVU9ZO1OJA8WA1wuok+gEb1Y9G1G/
TKeDj19oIEoWOsujlbm5/isEbfmS8yMQuE8rVVzMR5y3yz7F2nEDH1iUMXPwcxWx
wkIicpHGDr02mDMnWMe06zVB15sqXgCWtwYnepqsyhfpKyDmsTqhcn1XQg3Glzct
ufnvjPbHc3jK9GyyP99hyygjuVvBO2FmNvfxk1LSrhY=
`protect END_PROTECTED
