`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nUS7UsNNZBEfTkSUsCwQPTEmQSL/nIYtWnzOO2NwjLzabUJzctb9jn78+gB2SY6A
3PIYSbAj3iufcxGdxKggXBnXIfBROCUyvALshQ47299b7h0Ojo8Ki8HSueToOn34
5pGHLBrU8399IflGCeUlRpSVW30IGJvlLMdk56Mw9KN8hHw1/9LhSHwH2wiR7gGB
0WmWiLp1J28X+NFr4U+6w+1CcutibFeF9M4PWc36An3IRPN+RkCydmQH4xXZsaIP
gvI6oDK2kSYwRQDybwXZIoKi3BanzbQZn4QTr8oGFIXP8Uzy7OGsjgI8ITdvOray
4iUqzQ8iVA4f8ZEo97ebPjkH9HwZ81YwIG/8H9dGDmkwNZ+H//Y7vN1iOi/ryQ0u
tRvLV6rTXET0XRf4f4FjqwGfLwx4+Q6bxrygKBmlnumd2FTN7AkuRuFQ8VF9eUCI
alVJBmo0TSDN3KgEcns/vozVYCPvusiVlFpeW7Jq7xw12XUytWfk2GpDI/jsrUDn
Gn+dLvyYY8Y0HJBap7G3WX5tkFJIdeoJqz7US584d5AV1cyFUZumx94V6WIZVRvY
jkMA+ZJ8R8ucevP2PfmleM4flLst72TsZK2IEgO/m8MRw+aiag4Ser4xA/S8Ns1a
gkZwKiBNtuV9PiGfjWUR0w==
`protect END_PROTECTED
