`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t6UfT1Y+O5ViOErqDw8qUzfeNqryfb0kUXtzNNVzwWeEbLSykbBG5RL/Do2FmYK5
Uk+wAF4Sb+dW6m+NTPHzezGf1BGkHc6i/6HiI5g863AdOP2/VNTU5U7gtY68Pweb
Np1bHT4j2xNev/1kaNf+snhQIpPu8mnX9B/zgWoeziOBcCugIxxV3Em0X+NjwS+I
UOHlIyRRPSM5hCme9UhrTruuePoVkfxDZrzdqJqmZXhTOjwXUhoWqzdZpTa+qXdC
77yeUsN8avM+tXf3oOazS7GhuXXNgIPcOA6szYpiUrrfXsVocZ7MZkeRJ08TI9Tv
Y653ZS8z2+H+jJmJx3LG2vmKTFnkp5FkBQNGGfrO/xX5L+mgpL/q5lfULPkorg/X
bct6cRQD1xQ4E1taDmk4weYVpuUG1khxs7FdfvWfWgeQxaMUsUhn3NAgdsLyVOHN
Bti7PVlJRypbF8EHm8YFiex2zp2qGFcvqqrupvCBEqM1263RJv9sAEIRlsQybnX8
fZZt4YQVgMvTghyWhZT01Cr+YozwyQHKurXwK4+uU6A=
`protect END_PROTECTED
